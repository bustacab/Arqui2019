module imem #(parameter N = 32) (input logic  [5:0]   addr,
											output logic [N-1:0] q);

	
	logic [31:0] ROM [0:63] = '{32'hcb1e03de, 32'h8b040000, 32'h00000000, 32'h00000000, 
										32'h8b040001, 32'h00000000, 32'h00000000, 32'h8b040022, 
										32'h00000000, 32'h00000000, 32'h8b040043, 32'hf80003c0, 
										32'hf80083c1, 32'hf80103c2, 32'hf80183c3, 32'hb400001e, 
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
																				 
	
	always_comb
		q = ROM[addr];
	
endmodule


/* Ejercicio 1 Practico 2
32'hf8000000, 32'hf8008001, 32'hf8010002, 32'hf8018003,
										32'hf8020004, 32'hf8028005, 32'hf8030006, 32'hf8400007,
										32'hf8408008, 32'hf8410009, 32'hf841800a, 32'hf842000b,
										32'hf842800c, 32'hf843000d, 32'h00000000, 32'h00000000, 
										32'hcb0e01ce, 32'hb400004e, 32'hcb01000f, 32'h8b01000f, 
										32'h00000000, 32'h00000000, 32'hf803800f, 32'h00000000,
										32'h00000000, 32'h00000000, 32'hf803800f, 32'h00000000,
										32'h00000000, 32'h00000000, 32'hf803800f, 32'h00000000,
										32'h00000000, 32'h00000000, 32'hf803800f, 32'h00000000,
										32'h00000000, 32'h00000000, 32'hf803800f, 32'h00000000,
										32'h00000000, 32'h00000000, 32'hf803800f, 32'h00000000,
										32'h00000000, 32'h00000000, 32'hf803800f, 32'h00000000,
										32'h00000000, 32'h00000000, 32'hf803800f, 32'h00000000,
										32'h00000000, 32'h00000000, 32'hf803800f, 32'h00000000,
										32'h00000000, 32'h00000000, 32'hf803800f, 32'h00000000,
										32'h00000000, 32'h00000000, 32'hf803800f, 32'h00000000};

*/







/* Ejercicio 2 Lab

{32'hcb00001e, 32'h8b040001, 32'h00000000, 32'h00000000,
										32'h8b040022, 32'h00000000, 32'h00000000, 32'h8b040043,
										32'h00000000, 32'h00000000, 32'h8b040065, 32'hf80003c1,
										32'hf80083c2, 32'hf80103c3, 32'hf80183c5, 32'hb400001e,
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000,
										32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000};
*/
