module imem #(parameter N = 32) (input logic  [5:0]   addr,
											output logic [N-1:0] q);

	
	//logic [31:0] ROM [0:63] = '{32'hf8000000,32'hf8008001,32'hf8010002, // 1
	//									 32'hf8018003,32'hf8020004,32'hf8028005, // 2
	//									 32'hf8030006,32'hf8400007,32'hf8408008, // 3
	//									 32'hf8410009,32'hf841800a,32'hf842000b, // 4
	//									 32'hf842800c,32'hf843000d,32'hcb0e01ce, // 5
	//									 32'h00000000,32'h00000000,32'hb400004e, // 6
	//									 32'hcb01000f,32'h8b01000f,32'h00000000, // 7
	//									 32'h00000000,32'hf803800f,32'h00000000, // 8
	//									 32'h00000000,32'h00000000,32'h00000000, // 9
	//									 32'h00000000,32'h00000000,32'h00000000, // 10
	//									 32'h00000000,32'h00000000,32'h00000000, // 11
	//									 32'h00000000,32'h00000000,32'h00000000, // 12
	//									 32'h00000000,32'h00000000,32'h00000000, // 13
	//									 32'h00000000,32'h00000000,32'h00000000, // 14
	//									 32'h00000000,32'h00000000,32'h00000000, // 15
	//									 32'h00000000,32'h00000000,32'h00000000, // 16
	//									 32'h00000000,32'h00000000,32'h00000000, // 17
	//									 32'h00000000,32'h00000000,32'h00000000, // 18
	//									 32'h00000000,32'h00000000,32'h00000000, // 19
	//									 32'h00000000,32'h00000000,32'h00000000, // 20
	//									 32'h00000000,32'h00000000,32'h00000000, // 21
	//									 32'h00000000};
										 
	
	logic [31:0] ROM [0:63] = '{32'h91003c0a,32'haa14018b,32'h8a14018c, // 1
										 32'h8b0a0000,32'hcb01014a,32'hf800000b, // 2
										 32'hf800800c,32'hb5ffff8a,32'hf8010000, // 3
										 32'h00000000,32'h00000000,32'h00000000, // 4
										 32'h00000000,32'h00000000,32'h00000000, // 5
										 32'h00000000,32'h00000000,32'h00000000, // 6
										 32'h00000000,32'h00000000,32'h00000000, // 7
										 32'h00000000,32'h00000000,32'h00000000, // 8
										 32'h00000000,32'h00000000,32'h00000000, // 9
										 32'h00000000,32'h00000000,32'h00000000, // 10
										 32'h00000000,32'h00000000,32'h00000000, // 11
										 32'h00000000,32'h00000000,32'h00000000, // 12
										 32'h00000000,32'h00000000,32'h00000000, // 13
										 32'h00000000,32'h00000000,32'h00000000, // 14
										 32'h00000000,32'h00000000,32'h00000000, // 15
										 32'h00000000,32'h00000000,32'h00000000, // 16
										 32'h00000000,32'h00000000,32'h00000000, // 17
										 32'h00000000,32'h00000000,32'h00000000, // 18
										 32'h00000000,32'h00000000,32'h00000000, // 19
										 32'h00000000,32'h00000000,32'h00000000, // 20
										 32'h00000000,32'h00000000,32'h00000000, // 21
										 32'h00000000};
	
	
	always_comb
		q = ROM[addr];
	
endmodule


/* Whit NOP
'{32'hf8000000,32'hf8008001,32'hf8010002, // 1
32'hf8018003,32'hf8020004,32'hf8028005, // 2
32'hf8030006,32'hf8400007,32'hf8408008, // 3
32'hf8410009,32'hf841800a,32'hf842000b, // 4
32'hf842800c,32'hf843000d,32'hcb0e01ce, // 5
32'h00000000,32'h00000000,32'hb400004e, // 6
32'hcb01000f,32'h8b01000f,32'h00000000, // 7
32'h00000000,32'hf803800f,32'h00000000, // 8
32'h00000000,32'h00000000,32'h00000000, // 9
32'h00000000,32'h00000000,32'h00000000, // 10
32'h00000000,32'h00000000,32'h00000000, // 11
32'h00000000,32'h00000000,32'h00000000, // 12
32'h00000000,32'h00000000,32'h00000000, // 13
32'h00000000,32'h00000000,32'h00000000, // 14
32'h00000000,32'h00000000,32'h00000000, // 15
32'h00000000,32'h00000000,32'h00000000, // 16
32'h00000000,32'h00000000,32'h00000000, // 17
32'h00000000,32'h00000000,32'h00000000, // 18
32'h00000000,32'h00000000,32'h00000000, // 19
32'h00000000,32'h00000000,32'h00000000, // 20
32'h00000000,32'h00000000,32'h00000000, // 21
32'h00000000};
*/