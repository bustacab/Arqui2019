module muxs (input logic  a, b, s,
				 output logic y);

	mux(a, b, s, y);


endmodule
